// `include "./Main.v"
module tb_matrix;

reg CLK;
reg reset;
// wire [31:0] start;
// reg [31:0] WriteInstruction;

    main dut(
        .CLK(CLK),
        .reset(reset)
        // .start(start)
        // .hardcode(hardcode),
        // .start(start)
        // .WriteInstruction(WriteInstruction)
    );

        always
        #1 CLK<=~CLK;
        initial
        #1650 $finish;
    
initial begin
  $dumpfile("matrixtb.vcd");
  $dumpvars(0,tb_matrix);
  $readmemb("testinstr.mem",dut.f.im.memory);
  $readmemb("data.mem",dut.m.dm.memory);
  CLK = 1'b1;
  reset = 1'b1;#5;
  reset = 1'b0;#5;
  // start = 32'b0;#10;//b01110001001100010000000000000000;#10;
  // pc
  // WriteInstruction = 32'b01110001001100010000000000000000;   #10; // lw s1 t1 0
  // WriteInstruction = 32'b01110001001100010000000000000000;   #10;// lw s1 t1 0
  // WriteInstruction = 32'b00000001011010011010100000100000;   #10;// add s3 s1 s2 MULTIPLY
  // WriteInstruction = 32'b00000001011110111011100000100000;   #10;// add s4 s3 s4
  // WriteInstruction = 32'b01110001001100010000000000000001;   #10;// lw s1 t1 1
  // WriteInstruction = 32'b01110001010100100000000000000011;   #10;// lw s2 t2 3
  // WriteInstruction = 32'b00000001011010011010100000100000;   #10;// add s3 s1 s2 MULTIPLY
  // WriteInstruction = 32'b00000001011110111011100000100000;   #10;// add s4 s3 s4
  // WriteInstruction = 32'b01110001001100010000000000000010;   #10;// lw s1 t1 2
  // WriteInstruction = 32'b01110001010100100000000000000110;   #10;// lw s2 t2 6
  // WriteInstruction = 32'b00000001011010011010100000100000;   #10; // add s3 s1 s2 MULTIPLY
  // WriteInstruction = 32'b00000001011110111011100000100000;   #10;// add s4 s3 s4
  // WriteInstruction = 32'b10000001011100110000000000000000;   #10;// store s4 t3
/*  WriteInstruction =
  WriteInstruction =
			      32'h4000 : memory[0] = 32'b01110001001100010000000000000000; // lw s1 t1 0
            32'h4001 : memory[1] = 32'b01110001010100100000000000000000; // lw s2 t2 0
            32'h4002 : memory[2] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
            32'h4003 : memory[3] = 32'b00000001011110111011100000100000; // add s4 s3 s4
            32'h4000 : memory[4] = 32'b01110001001100010000000000000001; // lw s1 t1 1
            32'h4001 : memory[5] = 32'b01110001010100100000000000000011; // lw s2 t2 3
						32'h4002 : memory[6] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
						32'h4003 : memory[7] = 32'b00000001011110111011100000100000; // add s4 s3 s4
						32'h4000 : memory[8] = 32'b01110001001100010000000000000010; // lw s1 t1 2
						32'h4001 : memory[9] = 32'b01110001010100100000000000000110; // lw s2 t2 6
					  32'h4002 : memory[10] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
						32'h4003 : memory[11] = 32'b00000001011110111011100000100000; // add s4 s3 s4
						32'h4004 : memory[12] = 32'b10000001011100110000000000000000; // store s4 t3
						// 32'h4005 : memory[13] = 32'b00100001011110111000000000010001; // addi t3 t3 1
						// 32'h4004 : memory[14] = 32'b10000001011100110000000000000000; // store s4 t3

			            32'h4000 : memory[13] = 32'b01110001001100010000000000000000; // lw s1 t1 0
						32'h4001 : memory[14] = 32'b01110001010100100000000000000001; // lw s2 t2 1
						32'h4002 : memory[15] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
						32'h4003 : memory[16] = 32'b00000001011110111011100000100000; // add s4 s3 s4
						32'h4000 : memory[17] = 32'b01110001001100010000000000000001; // lw s1 t1 1
						32'h4001 : memory[18] = 32'b01110001010100100000000000000100; // lw s2 t2 4
						32'h4002 : memory[19] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
						32'h4003 : memory[20] = 32'b00000001011110111011100000100000; // add s4 s3 s4
						32'h4000 : memory[21] = 32'b01110001001100010000000000000010; // lw s1 t1 2
						32'h4001 : memory[22] = 32'b01110001010100100000000000000111; // lw s2 t2 7
						32'h4002 : memory[23] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
						32'h4003 : memory[24] = 32'b00000001011110111011100000100000; // add s4 s3 s4
						32'h4004 : memory[25] = 32'b10000001011100110000000000000001; // store s4 t3+1
						// 32'h4005 : memory[26] = 32'b00100001011110111000000000010010; // addi t3 t3 2
						// 32'h4004 : memory[27] = 32'b10000001011100110000000000000000; // store s4 t3

			            32'h4000 : memory[26] = 32'b01110001001100010000000000000000; // lw s1 t1 0
						32'h4001 : memory[27] = 32'b01110001010100100000000000000010; // lw s2 t2 2
						32'h4002 : memory[28] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
						32'h4003 : memory[29] = 32'b00000001011110111011100000100000; // add s4 s3 s4
						32'h4000 : memory[30] = 32'b01110001001100010000000000000001; // lw s1 t1 1
						32'h4001 : memory[31] = 32'b01110001010100100000000000000101; // lw s2 t2 5
						32'h4002 : memory[32] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
						32'h4003 : memory[33] = 32'b00000001011110111011100000100000; // add s4 s3 s4
						32'h4000 : memory[34] = 32'b01110001001100010000000000000010; // lw s1 t1 2
						32'h4001 : memory[35] = 32'b01110001010100100000000000001000; // lw s2 t2 8
						32'h4002 : memory[36] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
						32'h4003 : memory[37] = 32'b00000001011110111011100000100000; // add s4 s3 s4
						32'h4004 : memory[38] = 32'b10000001011100110000000000000010; // store s4 t3 + 2
						// 32'h4005 : memory[39] = 32'b00100001011110111000000000010011; // addi t3 t3 3
						// 32'h4004 : memory[40] = 32'b10000001011100110000000000000000; // store s4 t3

			            32'h4000 : memory[0] = 32'b01110001001100010000000000000011; // lw s1 t1 3
						32'h4001 : memory[1] = 32'b01110001010100100000000000000000; // lw s2 t2 0
						32'h4002 : memory[2] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
						32'h4003 : memory[3] = 32'b00000001011110111011100000100000; // add s4 s3 s4
						32'h4000 : memory[0] = 32'b01110001001100010000000000000100; // lw s1 t1 4
						32'h4001 : memory[1] = 32'b01110001010100100000000000000011; // lw s2 t2 3
						32'h4002 : memory[2] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
						32'h4003 : memory[3] = 32'b00000001011110111011100000100000; // add s4 s3 s4
						32'h4000 : memory[0] = 32'b01110001001100010000000000000101; // lw s1 t1 5
						32'h4001 : memory[1] = 32'b01110001010100100000000000000110; // lw s2 t2 6
						32'h4002 : memory[2] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
						32'h4003 : memory[3] = 32'b00000001011110111011100000100000; // add s4 s3 s4
						32'h4004 : memory[4] = 32'b10000001011100110000000000000000; // store s4 t3 + 3
						// 32'h4005 : memory[5] = 32'b00100001011110111000000000010100; // addi t3 t3 4
						// 32'h4004 : memory[4] = 32'b10000001011100110000000000000000; // store s4 t3

			            32'h4000 : memory[0] = 32'b01110001001100010000000000000011; // lw s1 t1 3
						32'h4001 : memory[1] = 32'b01110001010100100000000000000001; // lw s2 t2 1
						32'h4002 : memory[2] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
						32'h4003 : memory[3] = 32'b00000001011110111011100000100100; // add s4 s3 s4
						32'h4000 : memory[0] = 32'b01110001001100010000000000000100; // lw s1 t1 4
						32'h4001 : memory[1] = 32'b01110001010100100000000000000011; // lw s2 t2 4
						32'h4002 : memory[2] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
						32'h4003 : memory[3] = 32'b00000001011110111011100000100000; // add s4 s3 s4
						32'h4000 : memory[0] = 32'b01110001001100010000000000000101; // lw s1 t1 5
						32'h4001 : memory[1] = 32'b01110001010100100000000000000111; // lw s2 t2 7
						32'h4002 : memory[2] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
						32'h4003 : memory[3] = 32'b00000001011110111011100000100000; // add s4 s3 s4
						32'h4004 : memory[4] = 32'b10000001011100110000000000000000; // store s4 t3 + 4
						32'h4005 : memory[5] = 32'b00100001011110111000000000010001; // addi t3 t3 5
						32'h4004 : memory[4] = 32'b10000001011100110000000000000000; // store s4 t3

			            32'h4000 : memory[0] = 32'b01110001001100010000000000000011; // lw s1 t1 3
						32'h4001 : memory[1] = 32'b01110001010100100000000000000010; // lw s2 t2 2
						32'h4002 : memory[2] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
						32'h4003 : memory[3] = 32'b00000001011110111011100000100000; // add s4 s3 s4
						32'h4000 : memory[0] = 32'b01110001001100010000000000000100; // lw s1 t1 4
						32'h4001 : memory[1] = 32'b01110001010100100000000000000101; // lw s2 t2 5
						32'h4002 : memory[2] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
						32'h4003 : memory[3] = 32'b00000001011110111011100000100000; // add s4 s3 s4
						32'h4000 : memory[0] = 32'b01110001001100010000000000000101; // lw s1 t1 5
						32'h4001 : memory[1] = 32'b01110001010100100000000000001000; // lw s2 t2 8
						32'h4002 : memory[2] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
						32'h4003 : memory[3] = 32'b00000001011110111011100000100000; // add s4 s3 s4
						32'h4004 : memory[4] = 32'b10000001011100110000000000000101; // store s4 t3 + 5
						32'h4005 : memory[5] = 32'b00100001011110111000000000000110; // addi t3 t3 6
						32'h4004 : memory[4] = 32'b10000001011100110000000000000000; // store s4 t3

			      32'h4000 : memory[0] = 32'b01110001001100010000000000000110; // lw s1 t1 6
						32'h4001 : memory[1] = 32'b01110001010100100000000000000000; // lw s2 t2 0
						32'h4002 : memory[2] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
						32'h4003 : memory[3] = 32'b00000001011110111011100000100000; // add s4 s3 s4
						32'h4000 : memory[0] = 32'b01110001001100010000000000000111; // lw s1 t1 7
						32'h4001 : memory[1] = 32'b01110001010100100000000000000011; // lw s2 t2 3
						32'h4002 : memory[2] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
						32'h4003 : memory[3] = 32'b00000001011110111011100000100000; // add s4 s3 s4
						32'h4000 : memory[0] = 32'b01110001001100010000000000001000; // lw s1 t1 8
						32'h4001 : memory[1] = 32'b01110001010100100000000000000110; // lw s2 t2 6
						32'h4002 : memory[2] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
						32'h4003 : memory[3] = 32'b00000001011110111011100000100000; // add s4 s3 s4
						32'h4004 : memory[4] = 32'b10000001011100110000000000000110; // store s4 t3 + 6
						32'h4005 : memory[5] = 32'b00100001011110111000000000000111; // addi t3 t3 7
						32'h4004 : memory[4] = 32'b10000001011100110000000000000000; // store s4 t3

			      32'h4000 : memory[0] = 32'b01110001001100010000000000000110; // lw s1 t1 6
						32'h4001 : memory[1] = 32'b01110001010100100000000000000001; // lw s2 t2 1
						32'h4002 : memory[2] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
						32'h4003 : memory[3] = 32'b00000001011110111011100000100000; // add s4 s3 s4
						32'h4000 : memory[0] = 32'b01110001001100010000000000000111; // lw s1 t1 7
						32'h4001 : memory[1] = 32'b01110001010100100000000000000100; // lw s2 t2 4
						32'h4002 : memory[2] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
						32'h4003 : memory[3] = 32'b00000001011110111011100000100000; // add s4 s3 s4
						32'h4000 : memory[0] = 32'b01110001001100010000000000001000; // lw s1 t1 8
						32'h4001 : memory[1] = 32'b01110001010100100000000000000111; // lw s2 t2 7
						32'h4002 : memory[2] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
						32'h4003 : memory[3] = 32'b00000001011110111011100000100000; // add s4 s3 s4
						32'h4004 : memory[4] = 32'b10000001011100110000000000000111; // store s4 t3 + 7
						32'h4005 : memory[5] = 32'b00100001011110111000000000001000; // addi t3 t3 8
						32'h4004 : memory[4] = 32'b10000001011100110000000000000000; // store s4 t3

			      32'h4000 : memory[0] = 32'b01110001001100010000000000000110; // lw s1 t1 6
						32'h4001 : memory[1] = 32'b01110001010100100000000000000010; // lw s2 t2 2
						32'h4002 : memory[2] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
						32'h4003 : memory[3] = 32'b00000001011110111011100000100000; // add s4 s3 s4
						32'h4000 : memory[0] = 32'b01110001001100010000000000000111; // lw s1 t1 7
						32'h4001 : memory[1] = 32'b01110001010100100000000000000101; // lw s2 t2 5
						32'h4002 : memory[2] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
						32'h4003 : memory[3] = 32'b00000001011110111011100000100000; // add s4 s3 s4
						32'h4000 : memory[0] = 32'b01110001001100010000000000001000; // lw s1 t1 8
						32'h4001 : memory[1] = 32'b01110001010100100000000000001000; // lw s2 t2 8
						32'h4002 : memory[2] = 32'b00000001011010011010100000100000; // add s3 s1 s2 MULTIPLY
						32'h4003 : memory[3] = 32'b00000001011110111011100000100000; // add s4 s3 s4
						32'h4004 : memory[4] = 32'b10000001011100110000000000001000; // store s4 t3 + 8
						32'h4005 : memory[5] = 32'b00100001011110111000000000010001; // addi t3 t3 1
						32'h4004 : memory[4] = 32'b10000001011100110000000000000000; // store s4 t3
*/
end
endmodule
